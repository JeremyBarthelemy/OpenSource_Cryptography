
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
 
ENTITY ks_tb IS
END ks_tb;
 
ARCHITECTURE behavior OF ks_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT KoggeStone
    PORT(
         CLOCK : IN  std_logic;
         X : IN  std_logic_vector(255 downto 0);
         Y : IN  std_logic_vector(255 downto 0);
         S : OUT  std_logic_vector(255 downto 0);
         MUX_SEL : IN  std_logic;
         Save_Pin : IN  std_logic;
         Cin : IN  std_logic;
         Cout : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal CLOCK : std_logic := '0';
   signal X : std_logic_vector(255 downto 0) := (others => '0');
   signal Y : std_logic_vector(255 downto 0) := (others => '0');
   signal MUX_SEL : std_logic := '0';
   signal Save_Pin : std_logic := '0';
   signal Cin : std_logic := '0';

 	--Outputs
   signal S : std_logic_vector(255 downto 0);
   signal Cout : std_logic;

   -- Clock period definitions
   constant CLOCK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: KoggeStone PORT MAP (
          CLOCK => CLOCK,
          X => X,
          Y => Y,
          S => S,
          MUX_SEL => MUX_SEL,
          Save_Pin => Save_Pin,
          Cin => Cin,
          Cout => Cout
        );

   -- Clock process definitions
   CLOCK_process :process
   begin
		CLOCK <= '0';
		wait for CLOCK_period/2;
		CLOCK <= '1';
		wait for CLOCK_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		Cin <= '0';
		Save_Pin <= '1';
		X <= "0000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010";
		Y <= "0000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111111111111111111111111111111111111111111111111111111111111111";
		WAIT FOR CLOCK_PERIOD;
		Save_Pin <= '0';
		X <= (OTHERS => '1');
		Y <= "0111111111010011111111111111110000011010101011111111100000100010000000000000000000000001111010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101111111111111111111111111111111111111111111111111111111111111111100";
		WAIT FOR CLOCK_PERIOD*7;
		Cin <= '1';
		X <= "0000000000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010";
		Y <= "0000000000000000000000000000000000000000000011010100101010100101010010000101010111101010100000101111111111111111111111100101010010101111101011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010";
		Save_Pin <= '1';
      WAIT;
   end process;

END;
