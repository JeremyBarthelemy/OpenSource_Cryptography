LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PISO IS
    PORT( 
				Clk : IN STD_LOGIC;
				Input : IN STD_LOGIC_VECTOR (255 DOWNTO 0);
				ENABLE : IN STD_LOGIC;
				RESET : IN STD_LOGIC;
            Output : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
				MUX_SEL : IN STD_LOGIC
			);
END PISO;

ARCHITECTURE piso_arch OF PISO IS
SIGNAL REG_2_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_3_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_4_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_5_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_6_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_7_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_8_IN : STD_LOGIC_VECTOR(31 DOWNTO 0);

SIGNAL REG_1_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_2_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_3_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_4_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_5_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_6_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_7_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG_8_OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

WITH MUX_SEL SELECT
REG_2_IN <= REG_1_OUT WHEN '1',
				Input(223 DOWNTO 192) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_3_IN <= REG_2_OUT WHEN '1',
				Input(191 DOWNTO 160) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_4_IN <= REG_3_OUT WHEN '1',
				Input(159 DOWNTO 128) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_5_IN <= REG_4_OUT WHEN '1',
				Input(127 DOWNTO 96) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_6_IN <= REG_5_OUT WHEN '1',
				Input(95 DOWNTO 64) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_7_IN <= REG_6_OUT WHEN '1',
				Input(63 DOWNTO 32) WHEN OTHERS;

WITH MUX_SEL SELECT
REG_8_IN <= REG_7_OUT WHEN '1',
				Input(31 DOWNTO 0) WHEN OTHERS;
				

REG_1 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>Input(255 DOWNTO 224), Q=> REG_1_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_2 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_2_IN, Q=>REG_2_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_3 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_3_IN, Q=>REG_3_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_4 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_4_IN, Q=>REG_4_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_5 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_5_IN, Q=>REG_5_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_6 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_6_IN, Q=>REG_6_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_7 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_7_IN, Q=>REG_7_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

REG_8 : ENTITY work.REG(reg_arch)
		  PORT MAP(D=>REG_8_IN, Q=>REG_8_OUT, ENABLE=>ENABLE, RESET=>RESET, Clock=>Clk);

Output <= REG_8_OUT;

END piso_arch;

