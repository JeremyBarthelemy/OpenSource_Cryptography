LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SIPO IS
    PORT( 
				Clk   : IN STD_LOGIC;
				ENABLE : IN STD_LOGIC;
				RESET : IN STD_LOGIC;
				Input : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
            Output : OUT STD_LOGIC_VECTOR (255 DOWNTO 0)
			);
END SIPO;

ARCHITECTURE sipo_arch OF SIPO IS
SIGNAL REG1OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG2OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG3OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG4OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG5OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG6OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG7OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);
SIGNAL REG8OUT : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN

Reg_1 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>Input,Q=>REG1OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_2 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG1OUT,Q=>REG2OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_3 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG2OUT,Q=>REG3OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_4 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG3OUT,Q=>REG4OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_5 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG4OUT,Q=>REG5OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_6 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG5OUT,Q=>REG6OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_7 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG6OUT,Q=>REG7OUT,ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Reg_8 : ENTITY work.REG2(reg2_arch)
		PORT MAP(D=>REG7OUT,Q=>REG8OUT, ENABLE=>ENABLE,RESET=>RESET,CLOCK=>Clk);

Output <= REG1OUT & REG2OUT & REG3OUT & REG4OUT & REG5OUT & REG6OUT & REG7OUT & REG8OUT;

END sipo_arch;
